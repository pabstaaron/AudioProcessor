`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:26:12 10/13/2016 
// Design Name: 
// Module Name:    IFFTConfigDriver 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IFFTConfigDriver(
    input [3:0] frameSize,
    output [23:0] tData,
    output tValid,
    input tReady,
	 input CLK
    );


endmodule
